library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package hil_simulation_pkg is

    constant calculation_delay : integer := 1199;

end package hil_simulation_pkg;
